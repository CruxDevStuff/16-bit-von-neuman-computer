module computer(output out_m);
    reg outM = 0;

    assign out_m = outM; 
endmodule
