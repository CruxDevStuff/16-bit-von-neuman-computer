module ALU (input [15:0] x, y, output reg[15:0] out, out2, input zx, nx, zy, ny, f, no, output zr, ng);
    reg [15:0] x_in; 
    reg [15:0] y_in; 

    always @(x or y) begin
        if (zx) begin
            x_in = {16{1'b0}}; 
            out = x_in; 
        end else begin
            x_in = x;  
            out = x_in; 
        end

        if (nx) begin 
            x_in = ~x_in; 
            out = x_in;
        end 

        if (zy == 1'b1) begin
            y_in = {16{1'b0}}; 
            out2 = y_in; 
        end else begin
            y_in = y;  
            out2 = y_in; 
        end

        if (ny) begin 
            y_in = ~y_in; 
            out2 = y_in;
        end 
    end
endmodule

module AND_N(input [15:0] x, y, output [15:0] out); 
    parameter N = 16; 
    genvar i; 

    generate
        for (i = 0; i < N; i= i+1) begin
            and(out[i], x[i], y[i]); 
        end
    endgenerate
endmodule

module FULL_ADDER(input a, b, c, output sum, carry);
    wire sum1, carry1; 
    wire sum2, carry2; 

    xor(sum1, a, b); 
    and(carry1, a, b); 

    xor(sum, sum1, c); 
    and(carry2, sum1, c); 

    or(carry, carry1, carry2); 
endmodule


module ADDER_N(input [15:0] x, y, output [15:0] out); 
    parameter N = 16; // define the adder bit length. can be externally overwridden to change the adder size.
    wire [N-1:0] carry_out, sum_out; 

    genvar i; 

    generate
        for (i = 0; i < N; i= i+1) begin
            if (i==0)
                FULL_ADDER full_adder(x[i], y[i], 1'b0, out[i], carry_out[i]); 
            else
                FULL_ADDER full_adder(x[i], y[i], carry_out[i-1], out[i], carry_out[i]); 
        end
    endgenerate

endmodule
