module NOT(output out_val, input in_val);
	nand(out_val, in_val, 1); 
endmodule


// Use NAND gate as the primitive gate to build the rest of the gates
// NOT
// AND
// OR
// XOR
