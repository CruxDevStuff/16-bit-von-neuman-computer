module NOT(output out_val, input in_val);
	nand(out_val, in_val, 1); 
endmodule
